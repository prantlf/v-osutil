module main

fn main() {
	eprintln('stderr')
}
